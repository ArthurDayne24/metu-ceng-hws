`timescale 1ns / 1ps
module Data_Subsystem(
output  [23:0] MemAddr,
input [31:0] fromMemData,
output  [31:0] toMemData,
output  [31:0] Instr,
output  ZE,
output  NG,
output  CY,
output  OV,
input [4:0] AddrA,
input [4:0] AddrB,
input [4:0] AddrC,
input [3:0] ALUop,
input WrC,
input WrPC,
input WrCR,
input WrIR,
input Mem_ALU,
input PC_RA,
input IR_RB,
input ALU_PC,
input ZE_SE,
input Sin_Sout,
input Clk,
input Reset
    );
	 
	 
/*  DO NOT EDIT THIS FILE   */

	 
	 wire [31:0] DataA, DataB, DataC;
	 wire [31:0] Ain  , Bin; 
	 wire [31:0] ALUdata;
	 wire [31:0] tMemData;
	 wire [3:0]  Cond, CRout;
	 wire [31:0] IRreg, IRext;
	 wire [23:0] PCout;


	assign ZE = CRout[0];  
	assign CY = CRout[1];
	assign NG = CRout[2];  
	assign OV = CRout[3];
	assign Instr = IRreg;

	ALU ALU1(Ain,Bin,ALUop,ALUdata,Cond); 
	Reg_File GPR(AddrA,AddrB,AddrC,DataA,DataB,DataC,WrC,Reset,Clk);
	Register24 PC(ALUdata[23:0],PCout,WrPC,Reset,Clk);
	Register4 CR(Cond,CRout,WrCR,Reset,Clk);
	Register32 IR(tMemData,IRreg,WrIR,Reset,Clk);
	Mux32 MX1(tMemData,ALUdata,Mem_ALU,DataC);
	Mux32 MX2({8'b00000000,PCout},DataA,PC_RA,Ain);
	Extender ZSE(IRreg,ZE_SE,IRext);
	Mux32 MX3(IRext,DataB,IR_RB,Bin);
	Mux24 MX4(ALUdata[23:0],PCout,ALU_PC,MemAddr);
	Switch32 SL(fromMemData,toMemData,tMemData,DataB,Sin_Sout);



endmodule
